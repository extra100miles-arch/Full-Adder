library verilog;
use verilog.vl_types.all;
entity Test_sv_unit is
end Test_sv_unit;
