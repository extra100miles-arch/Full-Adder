library verilog;
use verilog.vl_types.all;
entity add_intf is
end add_intf;
