library verilog;
use verilog.vl_types.all;
entity Agent_sv_unit is
end Agent_sv_unit;
