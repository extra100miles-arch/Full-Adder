interface add_intf;
logic a;
logic b;
logic cin;
logic cout;
logic sum;
endinterface