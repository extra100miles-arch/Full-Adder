library verilog;
use verilog.vl_types.all;
entity my_package_sv_unit is
end my_package_sv_unit;
