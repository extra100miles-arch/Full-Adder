`include "uvm_macros.svh"
import uvm_pkg::*;
package my_package;
`include "Transaction.sv"
`include "Generator.sv"
`include "Driver.sv"
`include "Monitor.sv"
`include "Scoreboard.sv"
`include "Agent.sv"
`include "Environment.sv"
`include "Test.sv"
endpackage