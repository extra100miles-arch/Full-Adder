library verilog;
use verilog.vl_types.all;
entity my_packages is
end my_packages;
