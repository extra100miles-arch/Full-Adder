library verilog;
use verilog.vl_types.all;
entity Transaction_sv_unit is
end Transaction_sv_unit;
